--------------------------------------------------------------------------------
-- VHDL Architecture NSK600_lib.ram_s1.rtl
-- -----------------------------------------------------------------------------
-- Copyright (c) ABB Switzerland Ltd 2007
-- -----------------------------------------------------------------------------
-- Project      : O4CV
-- Library      : NSK600_lib
-- Unit         : ram_s1
-- Language     : VHDL
--------------------------------------------------------------------------------
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 74)
--
--------------------------------------------------------------------------------
-- $Workfile: ram_s1_rtl.vhd $
-- History:
-- $Log: /FPGA/NSK_FPGA/NSK600_lib/hdl_vm/ram_s1_rtl.vhd $ 
-- 
-- 9     11-07-06 9:40 Chstrue
-- R4 implementation
-- 
-- 6     07-10-11 15:23 Chmaglo1
-- -- no description --
-- 
-- 1     07-04-10 19:43 Chmaglo1
-- Variante: TDM Short Loop
-- 0     2007-04-02 13:37:10 Mathias Gloor (CH-L-0012267)
-- File Generated 
--
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
LIBRARY NSK600_lib;
USE NSK600_lib.typedef_p.all;

ENTITY ram_s1 IS
   PORT( 
      clk     : IN     std_logic;
      din     : IN     std_logic;
      rd_ptr  : IN     integer RANGE 0 TO 16383;
      reset_n : IN     std_logic;
      wr      : IN     std_logic;
      wr_ptr  : IN     integer RANGE 0 TO 16383;
      dout    : OUT    std_logic
   );

-- Declarations

END ram_s1 ;

--
--------------------------------------------------------------------------------
architecture rtl of ram_s1 is

-----------------------------------------------------------
-- Last edited:
--   110630: no changes
  
--------------------------------------------------------------------------------
-- DECLARATIONS
--------------------------------------------------------------------------------
type t_ram is array (0 to 16383) of std_logic; 
--signal ram : t_ram := X"1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788_1122334455667788";
signal ram : t_ram := (others=>'0');
attribute block_ram : boolean;
attribute block_ram of ram : signal is true;
--
begin
--------------------------------------------------------------------------------
-- PROCESSES
--------------------------------------------------------------------------------
process (clk)
begin
  if clk'event and clk = '1' then
    if wr = '1' then
      ram(wr_ptr) <= din;
    end if;
    dout <= ram(rd_ptr);
    
  end if;
end process;
--------------------------------------------------------------------------------
-- CONCURRENT LOGIC
--------------------------------------------------------------------------------
-- 
--------------------------------------------------------------------------------
end architecture rtl;
