--------------------------------------------------------------------------
-- $Workfile: tb_config_p_110215.vhd $
-- Part of	    :	ETL600 / MUX600
-- Language    :	VHDL
-- Created by	 :	Alexander Gygax, PTUKT2
-- Remarks	    :  
-- Purpose	    : 
-- Copyright	  :	ABB Switzerland Ltd. 2004
---------------------------------------------------------------------------
--
-- $Log: /FPGA/NSK_FPGA/NSK600_tb/hdl_vm/tb_config_p_110215.vhd $
-- 
-- 1     11-07-06 9:24 Chstrue
-- R4 implementation
-- 
-- 49    08-04-22 16:24 Chstrue
-- -- no description --
-- 
-- 48    6.09.06 13:51 Chalgyg
-- V.11 external clock master is not supported anymore, unless DUT is in
-- MUX mode.
-- 
-- 47    8.02.06 12:42 Chalgyg
-- Some bugs removed.
-- 
-- 46    20.01.06 9:26 Chalgyg
-- G.703 interface integrated.
-- 
-- 45    10.01.06 9:05 Chalgyg
-- LAN interface is now supported.
-- 
-- 43    16.06.05 10:39 Chalgyg
-- TC25: V.11 port 1 pattern changed.
-- 
-- 42    25.04.05 13:05 Chalgyg
-- TC15 repaired.
-- 
-- 41    18.04.05 15:57 Chalgyg
-- V.24 clock verify in TC10 to 12 disabled. Makes problems and no sense.
-- 
-- 40    14.04.05 13:21 Chalgyg
-- New Testcase added.
-- 
-- 39    13.04.05 10:39 Chalgyg
-- New TC added.
-- 
-- 38    7.04.05 16:28 Chalgyg
-- Added pattern_protocol.
-- 
-- 37    1.03.05 16:57 Chalgyg
-- -- no description --
-- 
-- 36    1.03.05 10:07 Chalgyg
-- Constant mux_sync_time added.
-- 
-- 35    24.02.05 15:10 Chalgyg
-- constant check_mux_frame added.
-- 
-- 33    10.02.05 15:47 Chalgyg
-- For DSP IF Test.
-- 
-- 32    7.02.05 11:49 Chalgyg
-- TC17 ... 20 changed.
-- 
-- 31    2.02.05 15:08 Chalgyg
-- 3 new testcases for V.11 check.
-- 
-- 30    24.01.05 13:28 Chalgyg
-- Frequency deviation limit for V.24 and V.11 port added.
-- 
-- 29    18.01.05 14:54 Chalgyg
-- -- no description --
-- 
-- 28    18.01.05 10:12 Chalgyg
-- mode_v11 added.
-- 
-- 27    23.12.04 11:57 Chalgyg
-- -- no description --
-- 
-- 26    23.12.04 11:14 Chalgyg
-- fs_jitter added.
-- 
-- 25    20.12.04 11:26 Chalgyg
-- start_delay added.
-- 
-- 24    17.12.04 13:18 Chalgyg
-- Delay check added.
-- 
-- 22    13.12.04 13:47 Chalgyg
-- -- no description --
-- 
-- 21    8.12.04 13:56 Chalgyg
-- Testcase 18 added.
-- 
-- 20    8.12.04 13:29 Chalgyg
-- -- no description --
-- 
-- 18    3.12.04 13:10 Chalgyg
-- -- no description --
-- 
-- 17    1.12.04 14:55 Chalgyg
-- Check_RXC added.
-- 
-- 15    22.10.04 16:24 Gygax02
-- -- no description --
-- 
-- 14    20.10.04 11:45 Gygax02
-- -- no description --
-- 
-- 12    14.10.04 16:23 Gygax02
-- -- no description --
-- 
-- 11    8.10.04 14:34 Gygax02
-- -- no description --
-- 
-- 10    7.10.04 17:10 Gygax02
-- -- no description --
-- 
-- 9     20.09.04 10:36 Unp00631
-- -- no description --
-- 
-- 8     19.08.04 11:05 Gygax02
-- -- no description --
-- 
---------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package tb_config_p is

  type t_modus is (reset,dsp_if_com,loop_fsk,out_adpsk,real_out,in_adpsk,loop_rts,loop_p_share,loop_v11,loop_mux_v11,loop_mux_v24,loop_mixed,loop_lan,loop_g703);
  subtype t_testcase is integer range 0 to 27;

  type testarray_int is array (0 to 5 , 0 to t_testcase'high) of integer;
  type testarray4_int is array (0 to 3 , 0 to t_testcase'high) of integer;
  type testarray_std_vec is array (0 to 5 , 0 to t_testcase'high) of std_logic_vector (7 downto 0);
  type testarray4_std_vec is array (0 to 3 , 0 to t_testcase'high) of std_logic_vector (7 downto 0);
  type tstarray11_std_vec7 is array (0 to 10 , 0 to t_testcase'high) of std_logic_vector (6 downto 0);
  type tstarray11_std_vec6 is array (0 to 10 , 0 to t_testcase'high) of std_logic_vector (5 downto 0);
  type testarray_std_log is array (0 to 3 , 0 to t_testcase'high) of std_logic;
  type testarray_char is array (0 to 5 , 0 to t_testcase'high) of character;
  type testvec_std_log is array (0 to t_testcase'high) of std_logic;
  type testvec_int is array (0 to t_testcase'high) of integer;
  type testvec_mod is array (0 to t_testcase'high) of t_modus;
  type testvec_char is array (0 to t_testcase'high) of character;
  type testvec_real is array (0 to t_testcase'high) of real;
  
  -- Comments                                                           |            |Sep. data in|     No flow|        Data|            |            |            |            |            |            |            |            |            |            |            |            |            |            |            | Inverted   | V.11 exter-|8bit pattern| FT1 pattern|   Incl. LAN|            |            |            |
  --                                                                    |            |RX/TX dir.  |     control|   sensitive|            |            |            |            |            |            |            |            |            |            |            |            |            |            |            |            | nal master |            |HW-Handshake| Incl. G.703|            |            |            |
  -- Testcase                                                     0            1            2            3            4            5            6            7            8            9          10           11           12           13           14           15           16           17           18           19           20           21           22           23           24           25           26           27
  constant dps_if_modus            : testvec_mod         :=  (     reset,  dsp_if_com,    loop_fsk,    loop_fsk,    loop_fsk,    loop_fsk,   out_adpsk,   out_adpsk,   out_adpsk,    real_out,    in_adpsk,    in_adpsk,    in_adpsk,    loop_rts,loop_p_share,loop_p_share,loop_p_share,    loop_v11,    loop_v11,    loop_v11,    loop_v11,loop_mux_v11,loop_mux_v24,loop_mux_v24,  loop_mixed,  loop_mixed,    loop_lan,   loop_g703); 

  constant do_testcase             : testvec_std_log     :=  (       '1',         '1',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '1',         '1',         '1',         '0');

  constant mode                    : testarray_char      := ((       'o',         'o',         'f',         'f',         'f',         'f',         'a',         'a',         'a',         'f',         'a',         'a',         'a',         'a',         's',         's',         's',         'o',         'o',         'o',         'o',         'o',         'm',         'm',         'm',         'm',         'o',         'o'),
                                                             (       'o',         'o',         'f',         'f',         'f',         'f',         'a',         'a',         'a',         'o',         'a',         'a',         'a',         'f',         's',         's',         'a',         'o',         'o',         'o',         'o',         'o',         'o',         'm',         'o',         'o',         'o',         'o'),
                                                             (       'o',         'o',         'f',         'f',         'f',         'f',         'a',         'a',         'a',         'o',         'a',         'a',         'a',         'a',         'o',         'o',         'a',         'o',         'o',         'o',         'o',         'o',         'o',         'm',         'o',         'o',         'o',         'o'),
                                                             (       'o',         'o',         'f',         'f',         'f',         'f',         'a',         'a',         'a',         'o',         'a',         'a',         'a',         'a',         'o',         'o',         'f',         'o',         'o',         'o',         'o',         'o',         'm',         'm',         'o',         'o',         'o',         'o'),
                                                             (       'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         's',         's',         's',         'o',         'o',         'o',         'o',         'o',         'o',         'm',         'o',         'o',         'o',         'o'),
                                                             (       'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         's',         's',         's',         'o',         'o',         'o',         'o',         'o',         'm',         'm',         'o',         'o',         'o',         'o'));
  
  constant switchbox_modem         : testvec_char        :=  (       'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'f',         'm',         'f',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o');

  constant baudrate_value_ofdm     : testvec_int         :=  (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,       14400,      307200,       64000,      128000,      256000,       28800,       56000,       12000,       96000,      320000,      320000,       56000,       72000);   -- in Bps

  constant baudrate_value          : testarray_int       := ((         0,           0,        1200,        1200,        4800,        2400,        9600,        4800,        2400,        9600,        2400,        4800,        2400,           0,        1200,        1200,        1200,           0,           0,           0,           0,           0,        2400,        2400,        1200,        1200,           0,           0),
                                                             (         0,           0,        2400,        1200,        9600,        4800,        4800,        2400,        9600,           0,        4800,        2400,        9600,           0,        1200,        1200,        2400,           0,           0,           0,           0,           0,           0,       19200,           0,           0,           0,           0),
                                                             (         0,           0,        4800,        1200,        1200,        9600,        2400,        9600,        4800,           0,        2400,        9600,        4800,           0,           0,           0,        9600,           0,           0,           0,           0,           0,           0,        1200,           0,           0,           0,           0),
                                                             (         0,           0,        9600,        1200,        2400,        1200,        2400,        4800,        9600,           0,        9600,        4800,        2400,           0,           0,           0,         600,           0,           0,           0,           0,           0,        2400,        2400,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,        1200,        1200,        1200,           0,           0,           0,           0,           0,           0,        9600,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,        1200,        1200,        1200,           0,           0,           0,           0,           0,        2400,        2400,           0,           0,           0,           0));  -- in Bps

  constant start_delay             : testvec_int         :=  (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0);   -- in us

  constant baudrate_deviation      : testarray_int       := ((         0,           0,          10,           0,        2000,         100,           0,           0,           0,           0,        -100,          10,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,        -500,           0,           0),
                                                             (         0,           0,         -20,           0,        4000,         200,           0,           0,           0,           0,         100,         -20,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,          50,           0,       -4000,        -200,           0,           0,           0,           0,         500,         300,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,         -30,           0,       -2000,        -100,           0,           0,           0,           0,        -500,           5,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0));  -- in ppm

  constant pattern_protocol        : testvec_char        :=  (       's',         's',         's',         's',         's',         's',         's',         's',         's',         's',         's',         's',         's',         's',         's',         's',         's',         's',         's',         's',         's',         's',         's',         'f',         's',         's',         's',         's');

  constant pattern_v24             : testarray_std_vec   := (("00000000",  "00000000",  "10111100",  "00100101",  "11001010",  "01101000",  "00000000",  "00000000",  "00000000",  "00000000",  "11001001",  "00000011",  "00111011",  "00000000",  "00000000",  "01111001",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "11100010",  "00000001",  "00110001",  "10101010",  "00000000",  "00000000"),
                                                             ("00000000",  "00000000",  "00100110",  "10101111",  "11001101",  "11101111",  "00000000",  "00000000",  "00000000",  "00000000",  "00000100",  "00010001",  "01000001",  "00000000",  "00000000",  "00000000",  "01100111",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000001",  "00000000",  "00000000",  "00000000",  "00000000"),
                                                             ("00000000",  "00000000",  "01011101",  "00001101",  "11111111",  "00001000",  "00000000",  "00000000",  "00000000",  "00000000",  "01101000",  "00000010",  "00110010",  "00000000",  "00000000",  "00000000",  "10111001",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000001",  "00000000",  "00000000",  "00000000",  "00000000"),
                                                             ("00000000",  "00000000",  "00010101",  "01100101",  "00000001",  "10000000",  "00000000",  "00000000",  "00000000",  "00000000",  "10000001",  "10000000",  "01000000",  "00000000",  "00000000",  "00000000",  "11110110",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "01110111",  "00000001",  "00000000",  "00000000",  "00000000",  "00000000"),
                                                             ("00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "01001101",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000001",  "00000000",  "00000000",  "00000000",  "00000000"),
                                                             ("00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "10111001",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00100100",  "00000001",  "00000000",  "00000000",  "00000000",  "00000000"));

  constant nr_of_repetitions_v24   : testarray_int       := ((         0,           0,           4,          16,          16,           8,           0,           0,           0,           0,           8,           8,           4,           0,           8,           8,           4,           0,           0,           0,           0,           0,           4,           1,          16,           4,           0,           0),
                                                             (         0,           0,           8,          16,          32,          16,           0,           0,           0,           0,          16,           4,          16,           0,           8,           8,           8,           0,           0,           0,           0,           0,           0,           1,           0,           0,           0,           0),
                                                             (         0,           0,          16,          16,           4,          32,           0,           0,           0,           0,           8,          16,           8,           0,           0,           0,          32,           0,           0,           0,           0,           0,           0,           1,           0,           0,           0,           0),
                                                             (         0,           0,          32,          16,           8,           4,           0,           0,           0,           0,          32,           8,           4,           0,           0,           0,           2,           0,           0,           0,           0,           0,           5,           1,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           8,           8,           4,           0,           0,           0,           0,           0,           0,           1,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           8,           8,           4,           0,           0,           0,           0,           0,           3,           1,           0,           0,           0,           0));
                                                           
  constant pattern_dsp_if          : testarray4_std_vec  := (("00000000",  "00000000",  "00110001",  "00000000",  "00000000",  "00000000",  "10101100",  "11101000",  "10100100",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000"),
                                                             ("00000000",  "00000000",  "11000110",  "00000000",  "00000000",  "00000000",  "00100101",  "10000000",  "11111101",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "01101001",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000"),
                                                             ("00000000",  "00000000",  "01010000",  "00000000",  "00000000",  "00000000",  "11101111",  "00001001",  "11101100",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000100",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000"),
                                                             ("00000000",  "00000000",  "00100111",  "00000000",  "00000000",  "00000000",  "10111100",  "10101100",  "00101000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000"));

  constant nr_of_repetitions_dsp   : testarray4_int      := ((         0,           0,           4,           0,           0,           0,          16,           8,           4,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           8,           0,           0,           0,           8,           4,          16,           0,           0,           0,           0,           0,           0,           0,           8,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,          16,           0,           0,           0,           4,          16,           8,           0,           0,           0,           0,           0,           0,           0,          32,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,          32,           0,           0,           0,           4,           8,          16,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0));

  constant jitter_amplitude        : testarray_int       := ((         0,           0,          20,           0,           0,          10,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,         100,           0,           0,         200,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           5,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           2,           0,           0,           5,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0));  -- in ns
                                                           
  constant jitter_frequency        : testarray_int       := ((         0,           0,         100,           0,           0,        1000,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,        2000,           0,           0,         500,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,          10,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,       10000,           0,           0,         800,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0));  -- in Hz
                                                           
  constant glitch_off_duration     : testarray_int       := ((         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0));  -- in us
                                                           
  constant glitch_on_duration      : testarray_int       := ((         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0));  -- in ps

  constant mode_v11                : testvec_char        :=  (       'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'o',         'm',         'o',         'o',         'o',         'o',         'm',         'o',         'o',         'm',         'm',         'm',         'm');

  constant baudrate_value_v11      : testarray4_int      := ((         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,       64000,       64000,      128000,      256000,       28800,        9600,           0,           0,        9600,       80000,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,      128000,           0,           0,           0,           0,       19200,           0,           0,           0,      144000,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,       64000),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,       48000,           0));  -- in bps

  constant baudrate_deviation_v11  : testarray4_int      := ((         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,         240,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,          92),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0));  -- in ppm

  constant pattern_v11             : testarray4_std_vec  := (("00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00101110",  "00101110",  "01100100",  "11000011",  "00011110",  "01110010",  "00000000",  "00000000",  "01010100",  "11101111",  "00000000",  "00000000"),
                                                             ("00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "01000011",  "00000000",  "00000000",  "00000000",  "00000000",  "10011100",  "00000000",  "00000000",  "00000000",  "00011010",  "00000000",  "00000000"),
                                                             ("00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "11010110"),
                                                             ("00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "00000000",  "01110010",  "00000000"));

  constant nr_of_repetitions_v11   : testarray4_int      := ((         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,          10,         500,         200,         200,          20,          40,           0,           0,         100,         334,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,          40,           0,           0,           0,           0,          80,           0,           0,           0,         600,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,         256),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,          32,           0));

  constant jitter_amplitude_v11    : testarray4_int      := ((         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0));  -- in ns
                                                           
  constant jitter_frequency_v11    : testarray4_int      := ((         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0));  -- in Hz

  constant glitch_off_duration_v11 : testarray4_int      := ((         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0));  -- in us
                                                           
  constant glitch_on_duration_v11  : testarray4_int      := ((         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0),
                                                             (         0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0,           0));  -- in ps

  constant port_config_registers   : tstarray11_std_vec7 := (( "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0010001",   "0010001",   "0010001",   "0010001",   "0010001",   "0000001",   "0010001",   "0010001",   "0010001",   "0010001",   "0010001",   "0010001",   "0010001"),   -- OFDM interface
                                                             ( "0000000",   "0000000",   "0000001",   "0010001",   "0000001",   "0000001",   "0000001",   "0000001",   "0000001",   "0000001",   "0000001",   "0000001",   "0000001",   "0000001",   "1000001",   "0000001",   "0000001",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000001",   "0000001",   "0000001",   "0000001",   "0000000",   "0000000"),   -- V.24 Port 1
                                                             ( "0000000",   "0000000",   "0000001",   "0010001",   "0000001",   "0000001",   "0000001",   "0000001",   "0000001",   "0000000",   "0000001",   "0000001",   "0000001",   "0000001",   "1000001",   "0000001",   "0000001",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000001",   "0000000",   "0000000",   "0000000",   "0000000"),   -- V.24 Port 2
                                                             ( "0000000",   "0000000",   "0000001",   "0000001",   "1000001",   "0000001",   "0000001",   "0000001",   "0000001",   "0000000",   "0000001",   "0000001",   "0000001",   "0000001",   "0000000",   "0000000",   "0000001",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000001",   "0000000",   "0000000",   "0000000",   "0000000"),   -- V.24 Port 3
                                                             ( "0000000",   "0000000",   "0000001",   "0000001",   "1000001",   "0000001",   "0000001",   "0000001",   "0000001",   "0000000",   "0000001",   "0000001",   "0000001",   "0000001",   "0000000",   "0000000",   "0000001",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000001",   "0000001",   "0000000",   "0000000",   "0000000",   "0000000"),   -- V.24 Port 4
                                                             ( "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "1000001",   "0000001",   "0000001",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000001",   "0000000",   "0000000",   "0000000",   "0000000"),   -- V.24 Port 5
                                                             ( "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "1000001",   "0000001",   "0000001",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000001",   "0000001",   "0000000",   "0000000",   "0000000",   "0000000"),   -- V.24 Port 6
                                                             ( "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0010001",   "0010001",   "0010001",   "0010001",   "0001001",   "0010001",   "0000000",   "0000000",   "0010001",   "0010001",   "0000000",   "0000000"),   -- V.11 Port 1
                                                             ( "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0010001",   "0000000",   "0000000",   "0000000",   "0000000",   "0010001",   "0000000",   "0000000",   "0000000",   "0010001",   "0000000",   "0000000"),   -- V.11 Port 2
                                                             ( "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0010001"),   -- G.703
                                                             ( "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0000000",   "0010001",   "0000000"));  -- LAN
  -- Bits 6 downto 0 (DAS,JAC,AON,LRC,LTR,TPT,POE)

  constant clock_config_registers  : tstarray11_std_vec6 := ((  "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000100",    "000100",    "000100",    "000100",    "000100",    "101100",    "000100",    "000100",    "000100",    "000100",    "000100",    "000100",    "000100"),   -- OFDM interface
                                                             (  "000000",    "000000",    "000010",    "000010",    "000010",    "000010",    "000110",    "000110",    "000110",    "000010",    "000110",    "000110",    "000110",    "000010",    "000010",    "000111",    "000010",    "000000",    "000000",    "000000",    "000000",    "000000",    "000111",    "000111",    "000111",    "000111",    "000000",    "000000"),   -- V.24 Port 1
                                                             (  "000000",    "000000",    "000010",    "000010",    "000010",    "000010",    "000110",    "000110",    "000110",    "000000",    "000110",    "000110",    "000110",    "000010",    "000010",    "000111",    "000110",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000111",    "000000",    "000000",    "000000",    "000000"),   -- V.24 Port 2
                                                             (  "000000",    "000000",    "000010",    "000010",    "000010",    "000010",    "000110",    "000110",    "000110",    "000000",    "000110",    "000110",    "000110",    "000010",    "000000",    "000000",    "000110",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000111",    "000000",    "000000",    "000000",    "000000"),   -- V.24 Port 3
                                                             (  "000000",    "000000",    "000010",    "000010",    "000010",    "000010",    "000110",    "000110",    "000110",    "000000",    "000110",    "000110",    "000110",    "000010",    "000000",    "000000",    "000010",    "000000",    "000000",    "000000",    "000000",    "000000",    "000111",    "000111",    "000000",    "000000",    "000000",    "000000"),   -- V.24 Port 4
                                                             (  "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000010",    "000111",    "000010",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000111",    "000000",    "000000",    "000000",    "000000"),   -- V.24 Port 5
                                                             (  "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000010",    "000111",    "000010",    "000000",    "000000",    "000000",    "000000",    "000000",    "000111",    "000111",    "000000",    "000000",    "000000",    "000000"),   -- V.24 Port 6
                                                             (  "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "001101",    "001101",    "001100",    "001100",    "101100",    "001100",    "000000",    "000000",    "001100",    "001101",    "000000",    "000000"),   -- V.11 Port 1
                                                             (  "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "001101",    "000000",    "000000",    "000000",    "000000",    "001101",    "000000",    "000000",    "000000",    "001101",    "000000",    "000000"),   -- V.11 Port 2
                                                             (  "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000101"),   -- G.703 
                                                             (  "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "000000",    "001100",    "000000"));  -- LAN
  -- Bits 6 downto 2 (IAC,ICT,ICP,RXC,ASY,CLR)
  constant ofdm_port_ber           : testvec_real        :=  (       0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0,         0.0);

  constant loop_data_on_dsp_if     : testvec_std_log     :=  (       '0',         '0',         '0',         '1',         '1',         '1',         '0',         '0',         '0',         '0',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1');
  constant check_regenerated_txd   : testvec_std_log     :=  (       '0',         '0',         '1',         '1',         '1',         '1',         '0',         '0',         '0',         '0',         '1',         '1',         '1',         '0',         '1',         '0',         '1',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0');
  constant check_regenerated_rxd   : testvec_std_log     :=  (       '0',         '0',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '0',         '0',         '0',         '0',         '0',         '1',         '1',         '1',         '0',         '0',         '0',         '0',         '0',         '1',         '1',         '1',         '1',         '0',         '0');
  constant check_rxc               : testvec_std_log     :=  (       '0',         '0',         '0',         '0',         '0',         '0',         '1',         '1',         '1',         '0',         '0',         '0',         '0',         '0',         '0',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1');
  constant check_signalling        : testvec_std_log     :=  (       '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '1',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0');
  constant check_delay             : testvec_std_log     :=  (       '0',         '0',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '0',         '0',         '0',         '0',         '0',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1',         '1');
  constant check_mux_frame         : testvec_std_log     :=  (       '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '0',         '1',         '1',         '0',         '0',         '0',         '0',         '1',         '1',         '1',         '0',         '1',         '1',         '0');

  constant dsp_waitstates          : integer             :=  2;
  constant max_v24_deviation       : integer             :=  700; -- in ppm
  constant max_v11_deviation       : integer             :=  700; -- in ppm
  constant max_g703_deviation      : integer             :=  100; -- in ppm
  constant fs_jitter               : time                :=  0 ns;
  constant mux_sync_time           : time                :=  20 ms;

  function baudrate2code(baudrate: integer) return std_logic_vector;
  function baudrate2config(baudrate: integer) return integer;
  function mode2code(mode: character; switchbox: character) return std_logic_vector;
  function v11_mode2code(v11_mode: character) return std_logic;
  function share2code(mode: character) return std_logic;
  function deviation2time(deviation: integer) return time;
    
end tb_config_p;
