--
-- VHDL Package Header NSK600_tb.real_data
--
-- Created:
--          by - CHALGYG.UNKNOWN (CH-W-2364)
--          at - 13:20:18 15.12.2004
--
-- using Mentor Graphics HDL Designer(TM) 2004.1 (Build 41)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
PACKAGE tb_real_data_p IS
-----------------------------------------------------------
-- Last edited:
--   110630: bug fix (of old bugs) and adapt to R4




  type t_rxd_vec is array (0 to 99) of std_logic_vector(7 downto 0);
  
  constant real_rxd: t_rxd_vec := ("00110110",
                                   "10000111",
                                   "10000111",
                                   "10000111",
                                   "11000000",
                                   "01010001",
                                   "01010001",
                                   "01010001",
                                   "11001010",
                                   "00111101",
                                   "10110110",
                                   "00011011",
                                   "01010110",
                                   "10000001",
                                   "10000001",
                                   "10110110",
                                   "01001010",
                                   "01001010",
                                   "01001010",
                                   "10111101",
                                   "00110110",
                                   "10011011",
                                   "11010101",
                                   "01001011",
                                   "11011110",
                                   "11011110",
                                   "11011110",
                                   "00111101",
                                   "00111101",
                                   "00111101",
                                   "10110110",
                                   "00011011",
                                   "01010110",
                                   "11001011",
                                   "01000001",
                                   "11010001",
                                   "11010001",
                                   "11010001",
                                   "00110110",
                                   "00110110",
                                   "00110110",
                                   "10011011",
                                   "11010101",
                                   "01001011",
                                   "11000000",
                                   "00110110",
                                   "11001010",
                                   "11001010",
                                   "11001010",
                                   "00011011",
                                   "00011011",
                                   "00011011",
                                   "01010110",
                                   "11001011",
                                   "01000001",
                                   "10110101",
                                   "01011110",
                                   "10111101",
                                   "10111101",
                                   "10111101",
                                   "00010101",
                                   "00010101",
                                   "00010101",
                                   "01001011",
                                   "11000000",
                                   "00110110",
                                   "11011110",
                                   "01010001",
                                   "10110110",
                                   "10110110",
                                   "10110110",
                                   "00000111",
                                   "00000111",
                                   "00000111",
                                   "01000001",
                                   "10110110",
                                   "01011110",
                                   "11010001",
                                   "01001010",
                                   "10011011",
                                   "10011011",
                                   "10011011",
                                   "11010110",
                                   "00000001",
                                   "00000001",
                                   "00110110",
                                   "11011110",
                                   "01010001",
                                   "11001010",
                                   "00111101",
                                   "10010101",
                                   "10010101",
                                   "10010101",
                                   "11001011",
                                   "01011110",
                                   "01011110",
                                   "01011110",
                                   "11010110",
                                   "01001011",
                                   "01001011");

  
END tb_real_data_p;
